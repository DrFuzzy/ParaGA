-------------------------------------------------------------------------------
-- Title      : ROM Package
-- Project    : GA
-------------------------------------------------------------------------------
-- File       : rom_pkg.vhd
-- Author     : George Doyamis & Kyriakos Deliparaschos (kdelip@mail.ntua.gr)
-- Company    : NTUA/IRAL
-- Created    : 14/09/2006
-- Last update: 20/11/06
-- Platform   : Modelsim, Synplify, ISE
-------------------------------------------------------------------------------
-- Description: This package holds the rom data of the numerous ROM's in the
--              design. Of course it cannot be parametrized
-------------------------------------------------------------------------------
-- Copyright (c) 2006 NTUA
-------------------------------------------------------------------------------
-- revisions  :
-- date        version  author  description
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- LIBRARIES
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.ga_pkg.all;

--------------------------------------------------------------------------------
-- PACKAGE DECLARATION
--------------------------------------------------------------------------------
package rom_pkg is

  ------------------------
  -- Coordinates Map 
  ------------------------
  constant resol : positive := 3;       -- townres
  constant towns : positive := 8;       -- num_towns

  subtype town_x_y is std_logic_vector(2*resol-1 downto 0);
  type    towns_x_y is array(0 to towns) of town_x_y;
  --                                         
  constant coord_rom : towns_x_y := towns_x_y'(

    "ZZZZZZ",
    "001001",
    "001010",
    "010100",
    "011101",
    "010000",
    "011011",
    "100001",
    "101011"



--"ZZZZZZZZZZZZZZZZ",
--"0000000100000001",
--"0000000100000010",
--"0000001000000100",
--"0000001100000101",
--"0000001000000000",
--"0000001100000011",
--"0000010000000001",
--"0000010100000011"


--"0000001100000110",
--"0000010000000111",
--"0000011000000111",
--"0000011100000110",
--"0000010100000101",
--"0000010100000100",
--"0000011000000010",
--"0000011100000001"

    );

  ------------------------
  -- Initial generation
  ------------------------
  constant pop_sz : positive := 8;
  subtype  init_gene is std_logic_vector(resol*(towns-1)-1 downto 0);
  type     init_genes is array(0 to pop_sz) of init_gene;
  --                                         
  constant init_gen_rom : init_genes := init_genes'(
-------------------------------------------------
-- Population Size = 8
-------------------------------------------------
-- Matlab init_genes8.mat
"ZZZZZZZZZZZZZZZZZZZZZ",
"001010111100011101110",
"010001111101110011100",
"100011110001010111101",
"010111100001101110011",
"001111100110011101010",
"011101001110111010100",
"011101100110111010001",
"001011101111100010110"
-------------------------------------------------
-- Population Size = 16
-------------------------------------------------
-- Matlab init_genes16.mat
--"ZZZZZZZZZZZZZZZZZZZZZ",
--"111011001101010100110",
--"111011110010101100001",
--"110001011101100010111",
--"110001111010100101011",
--"100111110101001010011",
--"001011101111010100110",
--"011111010110101001100",
--"111100101001010011110",
--"001111011010100110101",
--"110011100111001101010",
--"110101100111011010001",
--"101001011111110100010",
--"010100111011101110001",
--"101001100011111110010",
--"101010111110100011001",
--"100111001101011110010"
---------------------------------------------------
-- Population Size = 32
---------------------------------------------------
-- Matlab init_genes32.mat
--"ZZZZZZZZZZZZZZZZZZZZZ",
--"101011111110010001100",
--"001110111010100011101",
--"100110011101001111010",
--"011100101010111110001",
--"110001101111011100010",
--"110001101010111011100",
--"100011010111110001101",
--"001010110101100011111",
--"001101011100010111110",
--"011010101110001111100",
--"010101001100011110111",
--"101001100010111110011",
--"010011110001111100101",
--"110101100011111001010",
--"011100101111110010001",
--"011110001111101100010",
--"101110011111010001100",
--"101100111110010001011",
--"110001111011100010101",
--"010011110001100101111",
--"101111110010001100011",
--"001111011100010101110",
--"011110001111010101100",
--"111101010001100011110",
--"111001100010011110101",
--"100001110010011101111",
--"110010001100101111011",
--"001100010101111110011",
--"001010110111101100011",
--"010100101111011001110",
--"011010101111110001100",
--"010001110111100011101"
);
end package rom_pkg;


--------------------------------------------------------------------------------
-- PACKAGE BODY DECLARATION
--------------------------------------------------------------------------------


package body rom_pkg is
-- empty
end package body rom_pkg;
