-- empty test1.vhd file - 1.1 
